`timescale 100ns/1ns
module Bias_ReLU_simd #(
    parameter integer ARRAY_N = 16,
    parameter integer OUT_WIDTH = 32
)  (
    input wire  clk,
    input wire  reset,
    input wire [$clog2(ARRAY_N) : 0]        w_index,
    input wire [OUT_WIDTH -1 : 0]           w_data,
    input wire                              w_en,

    input wire [ARRAY_N * OUT_WIDTH -1 : 0] data_in,
    input wire [ARRAY_N * OUT_WIDTH -1 : 0] data_out
);

reg [OUT_WITDH -1 : 0] bias_values [ARRAY_N -1 : 0];

always @(posedge clk)
begin
    if(w_en == 'b1)
    begin
        bias_values[w_index] <= w_data;
    end
end

wire data_out_0[ARRAY_N*OUT_WIDTH -1 : 0]

genvar i;
generate
for(i=0; i<ARRAY_N; i=i+1)
begin: SIMD_LOOP
    data_out_0[ARRAY_N * (i+1)-1 : ARRAY_N * (i)] = data_in[ARRAY_N * (i+1)-1 : ARRAY_N * (i)] + bias_values[i]
    data_out = [ARRAY_N * (i+1)-1 : ARRAY_N * (i)] = data_out_0[ARRAY_N * (i+1)-1] == 'b0 ? data_out_0[ARRAY_N * (i+1)-1 : ARRAY_N * (i)] : 0
end
endgenerate

endmodule
